netcdf xeoCoordinates {
dimensions:
	N_Lines_FR = 1280 ;
	N_Cols_FR = 4865 ;
variables:
	double longitude(N_Lines_FR, N_Cols_FR) ;
		longitude:long_name = "DEM_corrected_longitude" ;
		longitude:units = "degrees_east" ;
		longitude:valid_min = -180.0 ;
		longitude:valid_max = 180.0 ;
	double latitude(N_Lines_FR, N_Cols_FR) ;
		latitude:long_name = "DEM_geodetic_corrected_latitude" ;
		latitude:units = "degrees_north" ;
		latitude:valid_min = -90.0 ;
		latitude:valid_max = 90.0 ;
	short altitude(N_Lines_FR, N_Cols_FR) ;
		altitude:long_name = "DEM_corrected_altitude" ;
		altitude:units = "m" ;
		altitude:valid_min = -1000s ;
		altitude:valid_max = 9000s ;

// global attributes:
		:netCDF_version = "netCDF-4" ;
		:Conventions = "CF-1.4" ;
		:product_name = "${PRODUCT_NAME}" ;
		:data_set_name = "geoCoordinates" ;
		:title = "OL_1_EFR OLCI Level 1b Full Resolution Product, Geolocation Data Set" ;
		:institution = "ESRIN" ;
		:source = "test" ;
		:history = "generic" ;
		:input_files = "tbd" ;
		:auxiliary_files = "none" ;
		:references = "none" ;
		:contact = "tbd" ;
		:validity_start = "20101217T120000.0" ;
		:validity_stop = "20101217T130000.0" ;
		:creation_date = "20101217T140000.0" ;
		:absolute_orbit_number = 1U ;
		:spatial_resolution = 290s, 270s ;
data:
    latitude = ${LAT} ;
    longitude = ${LON} ;
}
