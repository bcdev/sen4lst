netcdf xeodetic_ao {
dimensions:
	nj = 960 ;
    ni = 1580 ;
variables:
	double latitude(nj, ni) ;
		latitude:long_name = "Latitude of detector FOV centre of the earth\'s surface" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:valid_min = -90.0 ;
		latitude:valid_max = 90.0 ;
	double longitude(nj, ni) ;
		longitude:long_name = "Longitude of detector FOV centre the earth\'s surface" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:valid_min = -180.0 ;
		longitude:valid_max = 180.0 ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "Full resolution Cartesian coordinates Annotation Data Sets" ;
		:institution = "ESRIN" ;
		:source = "test" ;
		:history = "generic" ;
		:comment = "no comments" ;
		:references = "none" ;
		:contact = "tbd" ;
		:netCDF_version = "netCDF-4" ;
		:processor_version = "2.0" ;
		:dataset_version = "2.0" ;
		:package_name = "${PRODUCT_NAME}.SAFE" ;
		:dataset_name = "geodetic_ao.nc" ;
		:dataset_type = "Measurement_Data_Set" ;
		:creation_time = "20101217T140000.0" ;
		:start_time = "20101217T120000.0" ;
		:stop_time = "20101217T130000.0" ;
		:resolution = 500s ;
		:start_offset = 0. ;
		:track_offset = 0. ;
data:
    latitude = ${LAT} ;
    longitude = ${LON} ;
}
